netcdf delme2 {
dimensions:
	lev = 2 ;
	time = 3 ;
	lat = 3 ;
	lon = 4 ;
	nbnd = 2 ;
variables:
	double time(time) ;
		time:standard_name = "time" ;
		time:units = "days since 2018-12-01" ;
		time:calendar = "365_day" ;
		time:bounds = "time_bnds" ;
	double lev(lev) ;
		lev:computed_standard_name = "air_pressure" ;
		lev:standard_name = "atmosphere_sigma_coordinate" ;
		lev:formula_terms = "sigma: a ptop: ptop ps: ps" ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:bounds = "lat_bnds" ;
		lat:units = "degrees_north" ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:bounds = "lon_bnds" ;
		lon:units = "degrees_east" ;
	double lon_bnds(lon,nbnd) ;
	double lat_bnds(lat,nbnd) ;
	double time_bnds(time,nbnd) ;
	double a(lev) ;
                a:long_name = "Formula term a";
		a:units = "1" ;
	double ptop;
                ptop:standard_name = "air_pressure_at_top_of_atmosphere_model";
		ptop:units = "hPa" ;
	double ps(time,lat, lon) ;
		ps:standard_name = "surface_air_pressure" ;
		ps:units = "hPa" ;
	double ta(time,lev, lat, lon) ;
                ta:long_name = "Atmospheric Air Temperature" ;
		ta:cell_methods = "lat: longitude: mean time: mean" ;
		ta:project = "Samples" ;
		ta:units = "K" ;
		ta:standard_name = "air_temperature" ;

// global attributes:
	:Conventions = "CF-1.7" ;
data:

 time = 15.5, 45.5, 75.5 ;
 time_bnds = 1., 31., 31., 61., 61., 91. ;

 lev = .25, .75 ;

 lat = 10, 30, 50 ;
 lat_bnds = 0, 20, 20, 40, 40, 60 ;

 lon = 45., 135., 225., 315.;
 lon_bnds = 0., 90., 90., 180., 180., 270., 270., 360.;

 a = 0.25, .75 ;

 ptop = 20 ;

 ps =
  0, 1, 2, 3, 4, 5, 6, 7, 8,
  9, 10, 11, 12, 13, 14, 15, 16, 17 ;

 ta =
  0, 1, 2, 3, 4, 5, 6, 7, 8,
  9, 10, 11, 12, 13, 14, 15, 16, 17,
  18, 19, 20, 21, 22, 23, 24, 25, 26,
  27, 28, 29, 30, 31, 32, 33, 34, 35 ;
}
